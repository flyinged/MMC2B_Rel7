
library IEEE;
use IEEE.STD_LOGIC_1164.all;

package COMPONENTS is


COMPONENT AND2
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT AND2A
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT AND2B
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT AND3
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT AND3A
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT AND3B
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT AND3C
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT AO12
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT AO13
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT AO14
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT AO15
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT AO16
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT AO17
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT AO18
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT AO1
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT AO1A
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT AO1B
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT AO1C
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT AO1D
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT AO1E
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT AOI1
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT AOI1A
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT AOI1B
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT AOI1C
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT AOI1D
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT AOI5
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT AX1
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT AX1A
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT AX1B
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT AX1C
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT AX1D
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT AX1E
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT AXO1
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT AXO2
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT AXO3
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT AXO5
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT AXO6
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT AXO7
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT AXOI1
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT AXOI2
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT AXOI3
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT AXOI4
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT AXOI5
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT AXOI7
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT PLLINT 
    port(
               A         : in    STD_ULOGIC;
               Y         : out    STD_ULOGIC);
END COMPONENT;

COMPONENT BUFD
    port(
                A         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;

COMPONENT INVD
    port(
                A         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;

COMPONENT BIBUF
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
                Y                : out    STD_ULOGIC);
END COMPONENT;

COMPONENT BIBUF_MSS
    generic(
               ACT_PIN       : String  := "";
               ACT_CONFIG    : integer := 0 );  
  port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
                Y                : out    STD_ULOGIC);
END COMPONENT;

COMPONENT BIBUF_F_12
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BIBUF_F_12D
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BIBUF_F_12U
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BIBUF_F_16
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BIBUF_F_16D
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BIBUF_F_16U
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BIBUF_F_24
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BIBUF_F_24D
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BIBUF_F_24U
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BIBUF_F_8
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BIBUF_F_8D
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BIBUF_F_8U
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;

COMPONENT BIBUF_LVCMOS15
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BIBUF_LVCMOS15D
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BIBUF_LVCMOS15U
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BIBUF_LVCMOS18
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BIBUF_LVCMOS18D
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BIBUF_LVCMOS18U
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BIBUF_LVCMOS25
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BIBUF_LVCMOS25D
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BIBUF_LVCMOS25U
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BIBUF_LVCMOS33
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BIBUF_LVCMOS33D
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BIBUF_LVCMOS33U
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BIBUF_LVCMOS5
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BIBUF_LVCMOS5D
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BIBUF_LVCMOS5U
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BIBUF_PCI
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BIBUF_PCIX
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BIBUF_S_12
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BIBUF_S_12D
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BIBUF_S_12U
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BIBUF_S_16
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BIBUF_S_16D
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BIBUF_S_16U
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BIBUF_S_24
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BIBUF_S_24D
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BIBUF_S_24U
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BIBUF_S_8
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BIBUF_S_8D
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BIBUF_S_8U
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT CLKBUF
    port(
                PAD         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;

COMPONENT CLKBUF_LVCMOS15
    port(
                PAD         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT CLKBUF_LVCMOS18
    port(
                PAD         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT CLKBUF_LVCMOS25
    port(
                PAD         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT CLKBUF_LVCMOS33
    port(
                PAD         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT CLKBUF_LVCMOS5
    port(
                PAD         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT CLKBUF_LVDS
    port(
      PADP                           :  in    STD_ULOGIC;
      PADN                           :  in    STD_ULOGIC;
      Y                              :  out   STD_ULOGIC);
END COMPONENT;


COMPONENT CLKBUF_LVPECL
    port(
      PADP                           :  in    STD_ULOGIC;
      PADN                           :  in    STD_ULOGIC;
      Y                              :  out   STD_ULOGIC);
END COMPONENT;


COMPONENT CLKBUF_PCI
    port(
                PAD         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT CLKBUF_PCIX
    port(
                PAD         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT DFI0
   port(
	D     :   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	QN	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFI0C0
   port(
	D     :   in   STD_ULOGIC;
	CLR	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	QN	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFI0C1
   port(
	D     :   in   STD_ULOGIC;
	CLR	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	QN	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFI0E0
   port(
	D     :   in   STD_ULOGIC;
	E	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	QN	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFI0E0C0
   port(
	D     :   in   STD_ULOGIC;
	CLR	:   in   STD_ULOGIC;
	E	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	QN	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFI0E0C1
   port(
	D     :   in   STD_ULOGIC;
	CLR	:   in   STD_ULOGIC;
	E	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	QN	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFI0E0P0
   port(
	D     :   in   STD_ULOGIC;
	PRE	:   in   STD_ULOGIC;
	E	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	QN	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFI0E0P1
   port(
	D     :   in   STD_ULOGIC;
	PRE	:   in   STD_ULOGIC;
	E	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	QN	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFI0E1
   port(
	D     :   in   STD_ULOGIC;
	E	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	QN	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFI0E1C0
   port(
	D     :   in   STD_ULOGIC;
	CLR	:   in   STD_ULOGIC;
	E	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	QN	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFI0E1C1
   port(
	D     :   in   STD_ULOGIC;
	CLR	:   in   STD_ULOGIC;
	E	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	QN	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFI0E1P0
   port(
	D     :   in   STD_ULOGIC;
	PRE	:   in   STD_ULOGIC;
	E	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	QN	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFI0E1P1
   port(
	D     :   in   STD_ULOGIC;
	PRE	:   in   STD_ULOGIC;
	E	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	QN	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFI0P0
   port(
	D     :   in   STD_ULOGIC;
	PRE	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	QN	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFI0P1
   port(
	D     :   in   STD_ULOGIC;
	PRE	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	QN	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFI0P1C1
   port(
	D     :   in   STD_ULOGIC;
	PRE	:   in   STD_ULOGIC;
	CLR	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	QN	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFI1
   port(
	D     :   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	QN	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFI1C0
   port(
	D     :   in   STD_ULOGIC;
	CLR	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	QN	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFI1C1
   port(
	D     :   in   STD_ULOGIC;
	CLR	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	QN	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFI1E0
   port(
	D     :   in   STD_ULOGIC;
	E	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	QN	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFI1E0C0
   port(
	D     :   in   STD_ULOGIC;
	CLR	:   in   STD_ULOGIC;
	E	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	QN	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFI1E0C1
   port(
	D     :   in   STD_ULOGIC;
	CLR	:   in   STD_ULOGIC;
	E	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	QN	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFI1E0P0
   port(
	D     :   in   STD_ULOGIC;
	PRE	:   in   STD_ULOGIC;
	E	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	QN	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFI1E0P1
   port(
	D     :   in   STD_ULOGIC;
	PRE	:   in   STD_ULOGIC;
	E	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	QN	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFI1E1
   port(
	D     :   in   STD_ULOGIC;
	E	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	QN	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFI1E1C0
   port(
	D     :   in   STD_ULOGIC;
	CLR	:   in   STD_ULOGIC;
	E	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	QN	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFI1E1C1
   port(
	D     :   in   STD_ULOGIC;
	CLR	:   in   STD_ULOGIC;
	E	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	QN	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFI1E1P0
   port(
	D     :   in   STD_ULOGIC;
	PRE	:   in   STD_ULOGIC;
	E	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	QN	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFI1E1P1
   port(
	D     :   in   STD_ULOGIC;
	PRE	:   in   STD_ULOGIC;
	E	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	QN	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFI1P0
   port(
	D     :   in   STD_ULOGIC;
	PRE	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	QN	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFI1P1
   port(
	D     :   in   STD_ULOGIC;
	PRE	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	QN	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFI1P1C1
   port(
	D     :   in   STD_ULOGIC;
	PRE	:   in   STD_ULOGIC;
	CLR	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	QN	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFN0
   port(
	D     :   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	Q	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFN0C0
   port(
	D     :   in   STD_ULOGIC;
	CLR	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	Q	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFN0C1
   port(
	D     :   in   STD_ULOGIC;
	CLR	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	Q	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFN0E0
   port(
	D     :   in   STD_ULOGIC;
	E	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	Q	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFN0E0C0
   port(
	D     :   in   STD_ULOGIC;
	CLR	:   in   STD_ULOGIC;
	E	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	Q	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFN0E0C1
   port(
	D     :   in   STD_ULOGIC;
	CLR	:   in   STD_ULOGIC;
	E	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	Q	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFN0E0P0
   port(
	D     :   in   STD_ULOGIC;
	PRE	:   in   STD_ULOGIC;
	E	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	Q	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFN0E0P1
   port(
	D     :   in   STD_ULOGIC;
	PRE	:   in   STD_ULOGIC;
	E	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	Q	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFN0E1
   port(
	D     :   in   STD_ULOGIC;
	E	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	Q	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFN0E1C0
   port(
	D     :   in   STD_ULOGIC;
	CLR	:   in   STD_ULOGIC;
	E	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	Q	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFN0E1C1
   port(
	D     :   in   STD_ULOGIC;
	CLR	:   in   STD_ULOGIC;
	E	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	Q	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFN0E1P0
   port(
	D     :   in   STD_ULOGIC;
	PRE	:   in   STD_ULOGIC;
	E	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	Q	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFN0E1P1
   port(
	D     :   in   STD_ULOGIC;
	PRE	:   in   STD_ULOGIC;
	E	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	Q	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFN0P0
   port(
	D     :   in   STD_ULOGIC;
	PRE	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	Q	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFN0P1
   port(
	D     :   in   STD_ULOGIC;
	PRE	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	Q	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFN0P1C1
   port(
	D     :   in   STD_ULOGIC;
	PRE	:   in   STD_ULOGIC;
	CLR	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	Q	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFN1
   port(
	D     :   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	Q	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFN1C0
   port(
	D     :   in   STD_ULOGIC;
	CLR	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	Q	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFN1C1
   port(
	D     :   in   STD_ULOGIC;
	CLR	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	Q	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFN1E0
   port(
	D     :   in   STD_ULOGIC;
	E	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	Q	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFN1E0C0
   port(
	D     :   in   STD_ULOGIC;
	CLR	:   in   STD_ULOGIC;
	E	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	Q	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFN1E0C1
   port(
	D     :   in   STD_ULOGIC;
	CLR	:   in   STD_ULOGIC;
	E	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	Q	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFN1E0P0
   port(
	D     :   in   STD_ULOGIC;
	PRE	:   in   STD_ULOGIC;
	E	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	Q	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFN1E0P1
   port(
	D     :   in   STD_ULOGIC;
	PRE	:   in   STD_ULOGIC;
	E	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	Q	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFN1E1
   port(
	D     :   in   STD_ULOGIC;
	E	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	Q	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFN1E1C0
   port(
	D     :   in   STD_ULOGIC;
	CLR	:   in   STD_ULOGIC;
	E	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	Q	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFN1E1C1
   port(
	D     :   in   STD_ULOGIC;
	CLR	:   in   STD_ULOGIC;
	E	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	Q	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFN1E1P0
   port(
	D     :   in   STD_ULOGIC;
	PRE	:   in   STD_ULOGIC;
	E	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	Q	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFN1E1P1
   port(
	D     :   in   STD_ULOGIC;
	PRE	:   in   STD_ULOGIC;
	E	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	Q	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFN1P0
   port(
	D     :   in   STD_ULOGIC;
	PRE	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	Q	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFN1P1
   port(
	D     :   in   STD_ULOGIC;
	PRE	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	Q	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DFN1P1C1
   port(
	D     :   in   STD_ULOGIC;
	PRE	:   in   STD_ULOGIC;
	CLR	:   in   STD_ULOGIC;
	CLK	:   in   STD_ULOGIC;
	Q	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DLI0
   port(
	D     :   in   STD_ULOGIC;
	G	:   in   STD_ULOGIC;
	QN	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DLI0C0
   port(
	D     :   in   STD_ULOGIC;
	CLR	:   in   STD_ULOGIC;
	G	:   in   STD_ULOGIC;
	QN	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DLI0C1
   port(
	D     :   in   STD_ULOGIC;
	CLR	:   in   STD_ULOGIC;
	G	:   in   STD_ULOGIC;
	QN	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DLI0P0
   port(
	D     :   in   STD_ULOGIC;
	PRE	:   in   STD_ULOGIC;
	G	:   in   STD_ULOGIC;
	QN	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DLI0P1
   port(
	D     :   in   STD_ULOGIC;
	PRE	:   in   STD_ULOGIC;
	G	:   in   STD_ULOGIC;
	QN	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DLI0P1C1
   port(
	D     :   in   STD_ULOGIC;
	PRE	:   in   STD_ULOGIC;
	CLR	:   in   STD_ULOGIC;
	G	:   in   STD_ULOGIC;
	QN	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DLI1
   port(
	D     :   in   STD_ULOGIC;
	G	:   in   STD_ULOGIC;
	QN	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DLI1C0
   port(
	D     :   in   STD_ULOGIC;
	CLR	:   in   STD_ULOGIC;
	G	:   in   STD_ULOGIC;
	QN	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DLI1C1
   port(
	D     :   in   STD_ULOGIC;
	CLR	:   in   STD_ULOGIC;
	G	:   in   STD_ULOGIC;
	QN	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DLI1P0
   port(
	D     :   in   STD_ULOGIC;
	PRE	:   in   STD_ULOGIC;
	G	:   in   STD_ULOGIC;
	QN	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DLI1P1
   port(
	D     :   in   STD_ULOGIC;
	PRE	:   in   STD_ULOGIC;
	G	:   in   STD_ULOGIC;
	QN	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DLI1P1C1
   port(
	D     :   in   STD_ULOGIC;
	PRE	:   in   STD_ULOGIC;
	CLR	:   in   STD_ULOGIC;
	G	:   in   STD_ULOGIC;
	QN	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DLN0
   port(
	D     :   in   STD_ULOGIC;
	G	:   in   STD_ULOGIC;
	Q	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DLN0C0
   port(
	D     :   in   STD_ULOGIC;
	CLR	:   in   STD_ULOGIC;
	G	:   in   STD_ULOGIC;
	Q	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DLN0C1
   port(
	D     :   in   STD_ULOGIC;
	CLR	:   in   STD_ULOGIC;
	G	:   in   STD_ULOGIC;
	Q	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DLN0P0
   port(
	D     :   in   STD_ULOGIC;
	PRE	:   in   STD_ULOGIC;
	G	:   in   STD_ULOGIC;
	Q	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DLN0P1
   port(
	D     :   in   STD_ULOGIC;
	PRE	:   in   STD_ULOGIC;
	G	:   in   STD_ULOGIC;
	Q	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DLN0P1C1
   port(
	D     :   in   STD_ULOGIC;
	PRE	:   in   STD_ULOGIC;
	CLR	:   in   STD_ULOGIC;
	G	:   in   STD_ULOGIC;
	Q	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DLN1
   port(
	D     :   in   STD_ULOGIC;
	G	:   in   STD_ULOGIC;
	Q	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DLN1C0
   port(
	D     :   in   STD_ULOGIC;
	CLR	:   in   STD_ULOGIC;
	G	:   in   STD_ULOGIC;
	Q	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DLN1C1
   port(
	D     :   in   STD_ULOGIC;
	CLR	:   in   STD_ULOGIC;
	G	:   in   STD_ULOGIC;
	Q	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DLN1P0
   port(
	D     :   in   STD_ULOGIC;
	PRE	:   in   STD_ULOGIC;
	G	:   in   STD_ULOGIC;
	Q	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DLN1P1
   port(
	D     :   in   STD_ULOGIC;
	PRE	:   in   STD_ULOGIC;
	G	:   in   STD_ULOGIC;
	Q	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT DLN1P1C1
   port(
	D     :   in   STD_ULOGIC;
	PRE	:   in   STD_ULOGIC;
	CLR	:   in   STD_ULOGIC;
	G	:   in   STD_ULOGIC;
	Q	:  out  STD_ULOGIC);
END COMPONENT;



COMPONENT GND
    port(
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT INBUF
    port(
                PAD         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;

COMPONENT INBUF_MSS
    generic(
               ACT_PIN       : String  := "";
               ACT_CONFIG    : integer := 0 );  
    port(
                PAD         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;

COMPONENT INBUF_MCCC
    generic(
               ACT_PIN       : String  := "";
               ACT_CONFIG    : integer := 0 );  
    port(
                PAD         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;

COMPONENT INBUF_A
    port(
                PAD         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT INBUF_DA
    port( 
                PAD         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT INBUF_LVCMOS15
    port(
                PAD         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT INBUF_LVCMOS15D
    port(
                PAD         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT INBUF_LVCMOS15U
    port(
                PAD         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT INBUF_LVCMOS18
    port(
                PAD         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT INBUF_LVCMOS18D
    port(
                PAD         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;

COMPONENT INBUF_LVCMOS18U
    port(
                PAD         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT INBUF_LVCMOS25
    port(
                PAD         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT INBUF_LVCMOS25D
    port(
                PAD         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT INBUF_LVCMOS25U
    port(
                PAD         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT INBUF_LVCMOS33
    port(
                PAD         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT INBUF_LVCMOS33D
    port(
                PAD         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT INBUF_LVCMOS33U
    port(
                PAD         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT INBUF_LVCMOS5
    port(
                PAD         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT INBUF_LVCMOS5D
    port(
                PAD         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;

COMPONENT INBUF_LVCMOS5U
    port(
                PAD         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT INBUF_LVDS
    port(
      PADP                           :  in    STD_ULOGIC;
      PADN                           :  in    STD_ULOGIC;
      Y                              :  out   STD_ULOGIC);

END COMPONENT;

COMPONENT INBUF_LVDS_MCCC
    generic(
               ACT_PIN       : String  := "");
    port(
      PADP                           :  in    STD_ULOGIC;
      PADN                           :  in    STD_ULOGIC;
      Y                              :  out   STD_ULOGIC);

END COMPONENT;

COMPONENT INBUF_LVPECL
    port(
      PADP                           :  in    STD_ULOGIC;
      PADN                           :  in    STD_ULOGIC;
      Y                              :  out   STD_ULOGIC);

END COMPONENT;

COMPONENT INBUF_LVPECL_MCCC
    generic(
               ACT_PIN       : String  := "");
  port(
      PADP                           :  in    STD_ULOGIC;
      PADN                           :  in    STD_ULOGIC;
      Y                              :  out   STD_ULOGIC);

END COMPONENT;

COMPONENT INBUF_PCI
    port(
                PAD         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT INBUF_PCIX
    port(
                PAD         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;

COMPONENT INV
    port(
                A         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;



COMPONENT MAJ3
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT MAJ3X
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT MAJ3XI
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT MIN3
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT MIN3X
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT MIN3XI
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT MX2
    port(
                A         : in    STD_ULOGIC;
                S         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT MX2A
    port(
                A         : in    STD_ULOGIC;
                S         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT MX2B
    port(
                A         : in    STD_ULOGIC;
                S         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT MX2C
    port(
                A         : in    STD_ULOGIC;
                S         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT NAND2
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT NAND2A
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT NAND2B
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;



COMPONENT NAND3
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT NAND3A
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT NAND3B
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT NAND3C
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT NOR2
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT NOR2A
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT NOR2B
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT NOR3
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT NOR3A
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT NOR3B
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT NOR3C
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT OA1
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT OA1A
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT OA1B
    port(
                C         : in    STD_ULOGIC;
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT OA1C
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT OAI1
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT OR2
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT OR2A
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT OR2B
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT OR3
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT OR3A
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT OR3B
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT OR3C
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT OUTBUF
    port(
                D         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT OUTBUF_MSS
    generic(
               ACT_PIN       : String  := "";
               ACT_CONFIG    : integer := 0 );  
  port(
                D         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;

COMPONENT OUTBUF_A
    port(
                D         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT OUTBUF_F_12
    port(
                D         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT OUTBUF_F_16
    port(
                D         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT OUTBUF_F_24
    port(
                D         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT OUTBUF_F_8
    port(
                D         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT OUTBUF_LVCMOS15
    port(
                D         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT OUTBUF_LVCMOS18
    port(
                D         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT OUTBUF_LVCMOS25
    port(
                D         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT OUTBUF_LVCMOS33
    port(
                D         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT OUTBUF_LVCMOS5
    port(
                D         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT OUTBUF_LVDS
    port(
      PADP                           :  out    STD_ULOGIC;
      PADN                           :  out    STD_ULOGIC;
      D                              :  in   STD_ULOGIC);

END COMPONENT;


COMPONENT OUTBUF_LVPECL
    port(
      PADP                           :  out    STD_ULOGIC;
      PADN                           :  out   STD_ULOGIC;
      D                              :  in   STD_ULOGIC);

END COMPONENT;


COMPONENT OUTBUF_PCI
    port(
                D         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT OUTBUF_PCIX
    port(
                D         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT OUTBUF_S_12
    port(
                D         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT OUTBUF_S_16
    port(
                D         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT OUTBUF_S_24
    port(
                D         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT OUTBUF_S_8
    port(
                D         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;

COMPONENT TRIBUFF_MSS
    generic(
               ACT_PIN       : String  := "";
               ACT_CONFIG    : integer := 0 );  
  port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;

COMPONENT TRIBUFF_F_12
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_F_12D
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_F_12U
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_F_16
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_F_16D
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_F_16U
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_F_24
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_F_24D
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_F_24U
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_F_8
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_F_8D
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_F_8U
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_LVCMOS15
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_LVCMOS15D
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_LVCMOS15U
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_LVCMOS18
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_LVCMOS18D
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_LVCMOS18U
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_LVCMOS25
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_LVCMOS25D
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_LVCMOS25U
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_LVCMOS33
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_LVCMOS33D
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_LVCMOS33U
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_LVCMOS5
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_LVCMOS5D
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_LVCMOS5U
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_PCI
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_PCIX
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_S_12
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_S_12D
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_S_12U
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_S_16
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_S_16D
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_S_16U
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_S_24
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_S_24D
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_S_24U
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_S_8
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_S_8D
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_S_8U
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT VCC
    port(
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT XA1
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT XA1A
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT XA1B
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT XA1C
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT XAI1
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT XAI1A
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT XNOR2
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT XNOR3
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT XO1
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT XO1A
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT XOR2
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT XOR3
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT ZOR3
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT ZOR3I
    port(
                A         : in    STD_ULOGIC;
                B         : in    STD_ULOGIC;
                C         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BUFF
    port(
                A         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT CLKINT 
  port(
                A         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT DDR_REG 
  port(
                D           : in    STD_ULOGIC;
                CLK         : in    STD_ULOGIC;
                CLR         : in    STD_ULOGIC;
                QR          : out    STD_ULOGIC;
                QF          : out    STD_ULOGIC);
END COMPONENT;

COMPONENT DDR_OUT 
  port(
                DR           : in    STD_ULOGIC;
                DF           : in    STD_ULOGIC;
                CLK          : in    STD_ULOGIC;
                CLR          : in    STD_ULOGIC;
                Q            : out    STD_ULOGIC);
END COMPONENT;


COMPONENT RAM4K9

    generic(
               MEMORYFILE       : String  := "");

    port(
               ADDRA0		: in    STD_ULOGIC;
               ADDRA1		: in    STD_ULOGIC;
               ADDRA2		: in    STD_ULOGIC;
               ADDRA3		: in    STD_ULOGIC;
               ADDRA4		: in    STD_ULOGIC;
               ADDRA5		: in    STD_ULOGIC;
               ADDRA6		: in    STD_ULOGIC;
               ADDRA7		: in    STD_ULOGIC;
               ADDRA8		: in    STD_ULOGIC;
               ADDRA9		: in    STD_ULOGIC;
               ADDRA10		: in    STD_ULOGIC;
               ADDRA11		: in    STD_ULOGIC;
               DINA0		: in    STD_ULOGIC;
               DINA1		: in    STD_ULOGIC;
               DINA2		: in    STD_ULOGIC;
               DINA3		: in    STD_ULOGIC;
               DINA4		: in    STD_ULOGIC;
               DINA5		: in    STD_ULOGIC;
               DINA6		: in    STD_ULOGIC;
               DINA7		: in    STD_ULOGIC;
               DINA8		: in    STD_ULOGIC;
               WIDTHA0		: in    STD_ULOGIC;
               WIDTHA1		: in    STD_ULOGIC;
               PIPEA		: in    STD_ULOGIC;
               WMODEA		: in    STD_ULOGIC;
               BLKA		: in    STD_ULOGIC;
               WENA		: in    STD_ULOGIC;
               CLKA		: in    STD_ULOGIC;
               ADDRB0           : in    STD_ULOGIC;
               ADDRB1           : in    STD_ULOGIC;
               ADDRB2           : in    STD_ULOGIC;
               ADDRB3           : in    STD_ULOGIC;
               ADDRB4           : in    STD_ULOGIC;
               ADDRB5           : in    STD_ULOGIC;
               ADDRB6           : in    STD_ULOGIC;
               ADDRB7           : in    STD_ULOGIC;
               ADDRB8           : in    STD_ULOGIC;
               ADDRB9           : in    STD_ULOGIC;
               ADDRB10          : in    STD_ULOGIC;
               ADDRB11          : in    STD_ULOGIC;
               DINB0            : in    STD_ULOGIC;
               DINB1            : in    STD_ULOGIC;
               DINB2            : in    STD_ULOGIC;
               DINB3            : in    STD_ULOGIC;
               DINB4            : in    STD_ULOGIC;
               DINB5            : in    STD_ULOGIC;
               DINB6            : in    STD_ULOGIC;
               DINB7            : in    STD_ULOGIC;
               DINB8            : in    STD_ULOGIC;
               WIDTHB0          : in    STD_ULOGIC;
               WIDTHB1          : in    STD_ULOGIC;
               PIPEB            : in    STD_ULOGIC;
               WMODEB           : in    STD_ULOGIC;
               BLKB             : in    STD_ULOGIC;
               WENB             : in    STD_ULOGIC;
               CLKB             : in    STD_ULOGIC;
               RESET		: in    STD_ULOGIC;
               DOUTA0		: out   STD_ULOGIC;
               DOUTA1           : out   STD_ULOGIC;
               DOUTA2           : out   STD_ULOGIC;
               DOUTA3           : out   STD_ULOGIC;
               DOUTA4           : out   STD_ULOGIC;
               DOUTA5           : out   STD_ULOGIC;
               DOUTA6           : out   STD_ULOGIC;
               DOUTA7           : out   STD_ULOGIC;
               DOUTA8           : out   STD_ULOGIC;
               DOUTB0           : out   STD_ULOGIC;
               DOUTB1           : out   STD_ULOGIC;
               DOUTB2           : out   STD_ULOGIC;
               DOUTB3           : out   STD_ULOGIC;
               DOUTB4           : out   STD_ULOGIC;
               DOUTB5           : out   STD_ULOGIC;
               DOUTB6           : out   STD_ULOGIC;
               DOUTB7           : out   STD_ULOGIC;
               DOUTB8           : out   STD_ULOGIC);
END COMPONENT;

COMPONENT RAM512X18

    generic(
               MEMORYFILE       : String  := "");

    port(
               RADDR0		: in    STD_ULOGIC;
               RADDR1           : in    STD_ULOGIC;
               RADDR2           : in    STD_ULOGIC;
               RADDR3           : in    STD_ULOGIC;
               RADDR4           : in    STD_ULOGIC;
               RADDR5           : in    STD_ULOGIC;
               RADDR6           : in    STD_ULOGIC;
               RADDR7           : in    STD_ULOGIC;
               RADDR8           : in    STD_ULOGIC;
               RW1		: in    STD_ULOGIC;
               RW0              : in    STD_ULOGIC;
               PIPE		: in    STD_ULOGIC;
               REN		: in    STD_ULOGIC;
               RCLK		: in    STD_ULOGIC;
               WADDR0		: in    STD_ULOGIC;
               WADDR1           : in    STD_ULOGIC;
               WADDR2           : in    STD_ULOGIC;
               WADDR3           : in    STD_ULOGIC;
               WADDR4           : in    STD_ULOGIC;
               WADDR5           : in    STD_ULOGIC;
               WADDR6           : in    STD_ULOGIC;
               WADDR7           : in    STD_ULOGIC;
               WADDR8           : in    STD_ULOGIC;
               WD0		: in    STD_ULOGIC;
               WD1		: in    STD_ULOGIC;
               WD2		: in    STD_ULOGIC;
               WD3		: in    STD_ULOGIC;
               WD4		: in    STD_ULOGIC;
               WD5		: in    STD_ULOGIC;
               WD6		: in    STD_ULOGIC;
               WD7		: in    STD_ULOGIC;
               WD8		: in    STD_ULOGIC;
               WD9		: in    STD_ULOGIC;
               WD10		: in    STD_ULOGIC;
               WD11		: in    STD_ULOGIC;
               WD12		: in    STD_ULOGIC;
               WD13		: in    STD_ULOGIC;
               WD14		: in    STD_ULOGIC;
               WD15		: in    STD_ULOGIC;
               WD16		: in    STD_ULOGIC;
               WD17		: in    STD_ULOGIC;
               WW1		: in    STD_ULOGIC;
               WW0              : in    STD_ULOGIC;
               WEN		: in    STD_ULOGIC;
               WCLK		: in    STD_ULOGIC;
               RESET		: in    STD_ULOGIC;
               RD0		: out   STD_ULOGIC;
               RD1              : out   STD_ULOGIC;
               RD2              : out   STD_ULOGIC;
               RD3              : out   STD_ULOGIC;
               RD4              : out   STD_ULOGIC;
               RD5              : out   STD_ULOGIC;
               RD6              : out   STD_ULOGIC;
               RD7              : out   STD_ULOGIC;
               RD8              : out   STD_ULOGIC;
               RD9              : out   STD_ULOGIC;
               RD10              : out   STD_ULOGIC;
               RD11              : out   STD_ULOGIC;
               RD12              : out   STD_ULOGIC; 
               RD13              : out   STD_ULOGIC;
               RD14              : out   STD_ULOGIC;
               RD15              : out   STD_ULOGIC;
               RD16              : out   STD_ULOGIC;
               RD17              : out   STD_ULOGIC);
END COMPONENT;

-- Removed for SAR28921 since the FLEXRAMs are not supported in SmartFusion
-- COMPONENT FLEXRAM4K9

    -- generic(
               -- MEMORYFILE       : String  := "");

    -- port(
               -- ADDRA0		: in    STD_ULOGIC;
               -- ADDRA1		: in    STD_ULOGIC;
               -- ADDRA2		: in    STD_ULOGIC;
               -- ADDRA3		: in    STD_ULOGIC;
               -- ADDRA4		: in    STD_ULOGIC;
               -- ADDRA5		: in    STD_ULOGIC;
               -- ADDRA6		: in    STD_ULOGIC;
               -- ADDRA7		: in    STD_ULOGIC;
               -- ADDRA8		: in    STD_ULOGIC;
               -- ADDRA9		: in    STD_ULOGIC;
               -- ADDRA10		: in    STD_ULOGIC;
               -- ADDRA11		: in    STD_ULOGIC;
               -- DINA0		: in    STD_ULOGIC;
               -- DINA1		: in    STD_ULOGIC;
               -- DINA2		: in    STD_ULOGIC;
               -- DINA3		: in    STD_ULOGIC;
               -- DINA4		: in    STD_ULOGIC;
               -- DINA5		: in    STD_ULOGIC;
               -- DINA6		: in    STD_ULOGIC;
               -- DINA7		: in    STD_ULOGIC;
               -- DINA8		: in    STD_ULOGIC;
               -- WIDTHA0		: in    STD_ULOGIC;
               -- WIDTHA1		: in    STD_ULOGIC;
               -- PIPEA		: in    STD_ULOGIC;
               -- WMODEA		: in    STD_ULOGIC;
               -- BLKA		: in    STD_ULOGIC;
               -- WENA		: in    STD_ULOGIC;
               -- CLKA		: in    STD_ULOGIC;
               -- ADDRB0           : in    STD_ULOGIC;
               -- ADDRB1           : in    STD_ULOGIC;
               -- ADDRB2           : in    STD_ULOGIC;
               -- ADDRB3           : in    STD_ULOGIC;
               -- ADDRB4           : in    STD_ULOGIC;
               -- ADDRB5           : in    STD_ULOGIC;
               -- ADDRB6           : in    STD_ULOGIC;
               -- ADDRB7           : in    STD_ULOGIC;
               -- ADDRB8           : in    STD_ULOGIC;
               -- ADDRB9           : in    STD_ULOGIC;
               -- ADDRB10          : in    STD_ULOGIC;
               -- ADDRB11          : in    STD_ULOGIC;
               -- DINB0            : in    STD_ULOGIC;
               -- DINB1            : in    STD_ULOGIC;
               -- DINB2            : in    STD_ULOGIC;
               -- DINB3            : in    STD_ULOGIC;
               -- DINB4            : in    STD_ULOGIC;
               -- DINB5            : in    STD_ULOGIC;
               -- DINB6            : in    STD_ULOGIC;
               -- DINB7            : in    STD_ULOGIC;
               -- DINB8            : in    STD_ULOGIC;
               -- WIDTHB0          : in    STD_ULOGIC;
               -- WIDTHB1          : in    STD_ULOGIC;
               -- PIPEB            : in    STD_ULOGIC;
               -- WMODEB           : in    STD_ULOGIC;
               -- BLKB             : in    STD_ULOGIC;
               -- WENB             : in    STD_ULOGIC;
               -- CLKB             : in    STD_ULOGIC;
               -- RESET		: in    STD_ULOGIC;
               -- DOUTA0		: out   STD_ULOGIC;
               -- DOUTA1           : out   STD_ULOGIC;
               -- DOUTA2           : out   STD_ULOGIC;
               -- DOUTA3           : out   STD_ULOGIC;
               -- DOUTA4           : out   STD_ULOGIC;
               -- DOUTA5           : out   STD_ULOGIC;
               -- DOUTA6           : out   STD_ULOGIC;
               -- DOUTA7           : out   STD_ULOGIC;
               -- DOUTA8           : out   STD_ULOGIC;
               -- DOUTB0           : out   STD_ULOGIC;
               -- DOUTB1           : out   STD_ULOGIC;
               -- DOUTB2           : out   STD_ULOGIC;
               -- DOUTB3           : out   STD_ULOGIC;
               -- DOUTB4           : out   STD_ULOGIC;
               -- DOUTB5           : out   STD_ULOGIC;
               -- DOUTB6           : out   STD_ULOGIC;
               -- DOUTB7           : out   STD_ULOGIC;
               -- DOUTB8           : out   STD_ULOGIC);
-- END COMPONENT;

-- COMPONENT FLEXRAM512X18

    -- generic(
               -- MEMORYFILE       : String  := "");

    -- port(
               -- RADDR0		: in    STD_ULOGIC;
               -- RADDR1           : in    STD_ULOGIC;
               -- RADDR2           : in    STD_ULOGIC;
               -- RADDR3           : in    STD_ULOGIC;
               -- RADDR4           : in    STD_ULOGIC;
               -- RADDR5           : in    STD_ULOGIC;
               -- RADDR6           : in    STD_ULOGIC;
               -- RADDR7           : in    STD_ULOGIC;
               -- RADDR8           : in    STD_ULOGIC;
               -- RW1		: in    STD_ULOGIC;
               -- RW0              : in    STD_ULOGIC;
               -- PIPE		: in    STD_ULOGIC;
               -- REN		: in    STD_ULOGIC;
               -- RCLK		: in    STD_ULOGIC;
               -- WADDR0		: in    STD_ULOGIC;
               -- WADDR1           : in    STD_ULOGIC;
               -- WADDR2           : in    STD_ULOGIC;
               -- WADDR3           : in    STD_ULOGIC;
               -- WADDR4           : in    STD_ULOGIC;
               -- WADDR5           : in    STD_ULOGIC;
               -- WADDR6           : in    STD_ULOGIC;
               -- WADDR7           : in    STD_ULOGIC;
               -- WADDR8           : in    STD_ULOGIC;
               -- WD0		: in    STD_ULOGIC;
               -- WD1		: in    STD_ULOGIC;
               -- WD2		: in    STD_ULOGIC;
               -- WD3		: in    STD_ULOGIC;
               -- WD4		: in    STD_ULOGIC;
               -- WD5		: in    STD_ULOGIC;
               -- WD6		: in    STD_ULOGIC;
               -- WD7		: in    STD_ULOGIC;
               -- WD8		: in    STD_ULOGIC;
               -- WD9		: in    STD_ULOGIC;
               -- WD10		: in    STD_ULOGIC;
               -- WD11		: in    STD_ULOGIC;
               -- WD12		: in    STD_ULOGIC;
               -- WD13		: in    STD_ULOGIC;
               -- WD14		: in    STD_ULOGIC;
               -- WD15		: in    STD_ULOGIC;
               -- WD16		: in    STD_ULOGIC;
               -- WD17		: in    STD_ULOGIC;
               -- WW1		: in    STD_ULOGIC;
               -- WW0              : in    STD_ULOGIC;
               -- WEN		: in    STD_ULOGIC;
               -- WCLK		: in    STD_ULOGIC;
               -- RESET		: in    STD_ULOGIC;
               -- RD0		: out   STD_ULOGIC;
               -- RD1              : out   STD_ULOGIC;
               -- RD2              : out   STD_ULOGIC;
               -- RD3              : out   STD_ULOGIC;
               -- RD4              : out   STD_ULOGIC;
               -- RD5              : out   STD_ULOGIC;
               -- RD6              : out   STD_ULOGIC;
               -- RD7              : out   STD_ULOGIC;
               -- RD8              : out   STD_ULOGIC;
               -- RD9              : out   STD_ULOGIC;
               -- RD10              : out   STD_ULOGIC;
               -- RD11              : out   STD_ULOGIC;
               -- RD12              : out   STD_ULOGIC; 
               -- RD13              : out   STD_ULOGIC;
               -- RD14              : out   STD_ULOGIC;
               -- RD15              : out   STD_ULOGIC;
               -- RD16              : out   STD_ULOGIC;
               -- RD17              : out   STD_ULOGIC);
-- END COMPONENT;

COMPONENT FIFO4K18
         port(
              RW0		: in    STD_ULOGIC;
              RW1		: in    STD_ULOGIC;
              RW2		: in    STD_ULOGIC;
              WW0		: in    STD_ULOGIC;
              WW1		: in    STD_ULOGIC;
              WW2		: in    STD_ULOGIC;
              ESTOP		: in    STD_ULOGIC;
              FSTOP		: in    STD_ULOGIC;
              AEVAL11		: in    STD_ULOGIC;
              AEVAL10           : in    STD_ULOGIC;
              AEVAL9           : in    STD_ULOGIC; 
              AEVAL8		: in    STD_ULOGIC;
              AEVAL7		: in    STD_ULOGIC;
              AEVAL6		: in    STD_ULOGIC;
              AEVAL5		: in    STD_ULOGIC;
              AEVAL4		: in    STD_ULOGIC;
              AEVAL3		: in    STD_ULOGIC;
              AEVAL2		: in    STD_ULOGIC;
              AEVAL1		: in    STD_ULOGIC;
              AEVAL0		: in    STD_ULOGIC;
              AFVAL11           : in    STD_ULOGIC;
              AFVAL10           : in    STD_ULOGIC;
              AFVAL9           : in    STD_ULOGIC; 
              AFVAL8            : in    STD_ULOGIC;
              AFVAL7            : in    STD_ULOGIC;
              AFVAL6            : in    STD_ULOGIC;
              AFVAL5            : in    STD_ULOGIC;
              AFVAL4            : in    STD_ULOGIC;
              AFVAL3            : in    STD_ULOGIC;
              AFVAL2            : in    STD_ULOGIC;
              AFVAL1            : in    STD_ULOGIC;
              AFVAL0            : in    STD_ULOGIC;
              REN		: in    STD_ULOGIC;
              RBLK		: in    STD_ULOGIC;
              RCLK		: in    STD_ULOGIC;
              WD17		: in    STD_ULOGIC;
              WD16		: in    STD_ULOGIC;
              WD15		: in    STD_ULOGIC;
              WD14		: in    STD_ULOGIC;
              WD13		: in    STD_ULOGIC;
              WD12		: in    STD_ULOGIC;
              WD11		: in    STD_ULOGIC;
              WD10		: in    STD_ULOGIC;
              WD9		: in    STD_ULOGIC;
              WD8		: in    STD_ULOGIC;
              WD7		: in    STD_ULOGIC;
              WD6		: in    STD_ULOGIC;
              WD5		: in    STD_ULOGIC;
              WD4		: in    STD_ULOGIC;
              WD3		: in    STD_ULOGIC;
              WD2		: in    STD_ULOGIC;
              WD1		: in    STD_ULOGIC;
              WD0		: in    STD_ULOGIC;
              WEN		: in    STD_ULOGIC;
              WBLK		: in    STD_ULOGIC;
              WCLK		: in    STD_ULOGIC;
              RPIPE		: in    STD_ULOGIC;
              RESET		: in    STD_ULOGIC;
              RD0		: out   STD_ULOGIC;
              RD1		: out   STD_ULOGIC;
              RD2		: out   STD_ULOGIC;
              RD3		: out   STD_ULOGIC;
              RD4		: out   STD_ULOGIC;
              RD5		: out   STD_ULOGIC;
              RD6		: out   STD_ULOGIC;
              RD7		: out   STD_ULOGIC;
              RD8		: out   STD_ULOGIC;
              RD9		: out   STD_ULOGIC;
              RD10		: out   STD_ULOGIC;
              RD11		: out   STD_ULOGIC;
              RD12		: out   STD_ULOGIC;
              RD13		: out   STD_ULOGIC;
              RD14		: out   STD_ULOGIC;
              RD15		: out   STD_ULOGIC;
              RD16		: out   STD_ULOGIC;
              RD17		: out   STD_ULOGIC;
              FULL		: out   STD_ULOGIC;
              AFULL		: out   STD_ULOGIC;
              EMPTY		: out   STD_ULOGIC;
              AEMPTY		: out   STD_ULOGIC);
END COMPONENT; 		 
 


COMPONENT BIBUF_F_2
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BIBUF_F_2D
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BIBUF_F_2U
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BIBUF_F_4
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BIBUF_F_4D
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BIBUF_F_4U
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BIBUF_F_6
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BIBUF_F_6D
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BIBUF_F_6U
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BIBUF_S_2
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BIBUF_S_2D
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BIBUF_S_2U
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BIBUF_S_4
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BIBUF_S_4D
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BIBUF_S_4U
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BIBUF_S_6
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BIBUF_S_6D
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT BIBUF_S_6U
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT OUTBUF_F_2
    port(
                D         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT OUTBUF_F_4
    port(
                D         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT OUTBUF_F_6
    port(
                D         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT OUTBUF_S_2
    port(
                D         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT OUTBUF_S_4
    port(
                D         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT OUTBUF_S_6
    port(
                D         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;



COMPONENT TRIBUFF_F_2
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_F_2D
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_F_2U
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_F_4
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_F_4D
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_F_4U
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_F_6
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_F_6D
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_F_6U
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_S_2
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_S_2D
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_S_2U
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_S_4
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_S_4D
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_S_4U
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_S_6
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_S_6D
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT TRIBUFF_S_6U
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT CLKDLY
  port (
        CLK         : in    STD_ULOGIC;
        DLYGL0       : in    STD_ULOGIC;
        DLYGL1       : in    STD_ULOGIC;
        DLYGL2       : in    STD_ULOGIC;
        DLYGL3       : in    STD_ULOGIC;
        DLYGL4       : in    STD_ULOGIC;
        GL         :  out    STD_ULOGIC);
END COMPONENT;

COMPONENT UJTAG
  port
    (
      UIREG0 : out std_logic;
      UIREG1 : out std_logic;
      UIREG2 : out std_logic;
      UIREG3 : out std_logic;
      UIREG4 : out std_logic;
      UIREG5 : out std_logic;
      UIREG6 : out std_logic;
      UIREG7 : out std_logic;
      URSTB : out std_logic;
      UDRCK : out std_logic;
      UDRCAP : out std_logic;
      UDRSH : out std_logic;
      UDRUPD : out std_logic;
      UTDI : out std_logic;
      UTDO : in std_logic;
      TDO : out std_logic;
      TMS : in std_logic;
      TDI : in std_logic;
      TCK : in std_logic;
      TRSTB : in std_logic
    );
END COMPONENT;

COMPONENT CLKBIBUF
    port(
                D               : in    STD_ULOGIC;
                E               : in    STD_ULOGIC;
                PAD             : inout STD_ULOGIC;
                Y               : out    STD_ULOGIC);
END COMPONENT;


COMPONENT CLKSRC
  port(
               A                : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;


COMPONENT RCOSC 
    port (
         CLKOUT            : out   STD_ULOGIC 
         );
END COMPONENT;


COMPONENT BIBUF_LVDS
    port(
          D            : in    STD_ULOGIC;
          E            : in    STD_ULOGIC;
          PADP, PADN   : inout STD_ULOGIC;
          Y            : out   STD_ULOGIC);
END COMPONENT;

COMPONENT TRIBUFF_LVDS
    port(
          D            : in    STD_ULOGIC;
          E            : in    STD_ULOGIC;
          PADP, PADN   : out   STD_ULOGIC);
END COMPONENT;

COMPONENT SIMBUF
    PORT(
                D         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;

COMPONENT BIBUF_OPEND_MSS
    generic(
               ACT_PIN       : String  := "";
               ACT_CONFIG    : integer := 0 );    
    port(
                E         : in    STD_ULOGIC;
                PAD         : inout STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;

COMPONENT MSSINT
    port(
                A         : in    STD_ULOGIC;
               Y                : out    STD_ULOGIC);
END COMPONENT;

COMPONENT MSS_XTLOSC 
    port (
      XTL          : in STD_ULOGIC;
      CLKOUT            : out   STD_ULOGIC 
      );
END COMPONENT;

COMPONENT MSS_LPXTLOSC 
    port (
      LPXIN          : in STD_ULOGIC;
      CLKOUT            : out   STD_ULOGIC 
      );
END COMPONENT;

COMPONENT MSS_AHB 
  generic (
    ACT_CONFIG : integer := 0 ;
    ACT_FCLK   : integer  := 0 ;
    ACT_DIE   : string  := "" ;
    ACT_PKG   : string  := "");
   port (      
      MSSHADDR        : out std_logic_vector(19 downto 0);
      MSSHWDATA       : out std_logic_vector(31 downto 0);
      MSSHTRANS      : out std_logic_vector(1 downto 0);
      MSSHSIZE        : out std_logic_vector(1 downto 0);
      MSSHLOCK        : out std_logic;
      MSSHWRITE       : out std_logic;
      MSSHRDATA       : in std_logic_vector(31 downto 0);
      MSSHREADY       : in std_logic;
      MSSHRESP        : in std_logic;
      FABHADDR        : in std_logic_vector(31 downto 0);
      FABHWDATA       : in std_logic_vector(31 downto 0);
      FABHTRANS      : in std_logic_vector(1 downto 0);
      FABHSIZE        : in std_logic_vector(1 downto 0);
      FABHMASTLOCK    : in std_logic;
      FABHWRITE       : in std_logic;
      FABHSEL         : in std_logic;
      FABHREADY       : in std_logic;
      FABHRDATA       : out std_logic_vector(31 downto 0);
      FABHREADYOUT    : out std_logic;
      FABHRESP        : out std_logic;
      SYNCCLKFDBK     : in std_logic;
      CALIBOUT        : out std_logic;
      CALIBIN         : in std_logic;
      FABINT          : in std_logic;
      MSSINT          : out std_logic_vector(7 downto 0);
      WDINT           : out std_logic;
      F2MRESETn       : in std_logic;
      DMAREADY        : in std_logic_vector(1 downto 0);
      RXEV            : in std_logic;
      VRON            : in std_logic;
      M2FRESETn       : out std_logic;
      DEEPSLEEP       : out std_logic;
      SLEEP           : out std_logic;
      TXEV            : out std_logic;
      UART0CTSn       : in std_logic;
      UART0DSRn       : in std_logic;
      UART0RIn        : in std_logic;
      UART0DCDn       : in std_logic;
      UART0RTSn       : out std_logic;
      UART0DTRn       : out std_logic;
      UART1CTSn       : in std_logic;
      UART1DSRn       : in std_logic;
      UART1RIn        : in std_logic;
      UART1DCDn       : in std_logic;
      UART1RTSn       : out std_logic;
      UART1DTRn       : out std_logic;
      I2C0SMBUSNI     : in std_logic;
      I2C0SMBALERTNI  : in std_logic;
      I2C0BCLK        : in std_logic;
      I2C0SMBUSNO     : out std_logic;
      I2C0SMBALERTNO  : out std_logic;
      I2C1SMBUSNI     : in std_logic;
      I2C1SMBALERTNI  : in std_logic;
      I2C1BCLK        : in std_logic;
      I2C1SMBUSNO     : out std_logic;
      I2C1SMBALERTNO  : out std_logic;
      MACM2FTXD          : out std_logic_vector(1 downto 0);
      MACF2MRXD          : in std_logic_vector(1 downto 0);
      MACM2FTXEN         : out std_logic;
      MACF2MCRSDV        : in std_logic;
      MACF2MRXER         : in std_logic;
      MACF2MMDI          : in std_logic;
      MACM2FMDO          : out std_logic;
      MACM2FMDEN         : out std_logic;
      MACM2FMDC          : out std_logic;
      FABSDD0D        : in std_logic;
      FABSDD1D        : in std_logic;
      FABSDD2D        : in std_logic;
      FABSDD0CLK      : in std_logic;
      FABSDD1CLK      : in std_logic;
      FABSDD2CLK      : in std_logic;
      FABACETRIG      : in std_logic;
      ACEFLAGS  : out std_logic_vector(31 downto 0);
      CMP0            : out std_logic;
      CMP1            : out std_logic;
      CMP2            : out std_logic;
      CMP3            : out std_logic;
      CMP4            : out std_logic;
      CMP5            : out std_logic;
      CMP6            : out std_logic;
      CMP7            : out std_logic;
      CMP8            : out std_logic;
      CMP9            : out std_logic;
      CMP10           : out std_logic;
      CMP11           : out std_logic;
      LVTTL0EN      : in std_logic;
      LVTTL1EN      : in std_logic;
      LVTTL2EN      : in std_logic;
      LVTTL3EN      : in std_logic;
      LVTTL4EN      : in std_logic;
      LVTTL5EN      : in std_logic;
      LVTTL6EN      : in std_logic;
      LVTTL7EN      : in std_logic;
      LVTTL8EN      : in std_logic;
      LVTTL9EN      : in std_logic;
      LVTTL10EN     : in std_logic;
      LVTTL11EN     : in std_logic;
      LVTTL0        : out std_logic;
      LVTTL1        : out std_logic;
      LVTTL2        : out std_logic;
      LVTTL3        : out std_logic;
      LVTTL4        : out std_logic;
      LVTTL5        : out std_logic;
      LVTTL6        : out std_logic;
      LVTTL7        : out std_logic;
      LVTTL8        : out std_logic;
      LVTTL9        : out std_logic;
      LVTTL10       : out std_logic;
      LVTTL11       : out std_logic;
      PUFABn          : out std_logic;
      VCC15GOOD        : out std_logic;
      VCC33GOOD        : out std_logic;
      FCLK          : in std_logic;
      MACCLKCCC       : in std_logic;
      RCOSC           : in std_logic;
      MACCLK          : in std_logic;
      PLLLOCK         : in std_logic;
      MSSRESETn       : in std_logic;
      GPI             : in std_logic_vector(31 downto 0);
      GPO             : out std_logic_vector(31 downto 0);
      GPOE            : out std_logic_vector(31 downto 0);
      SPI0DO          : out std_logic;
      SPI0DOE         : out std_logic;
      SPI0DI          : in std_logic;
      SPI0CLKI        : in std_logic;
      SPI0CLKO        : out std_logic;
      SPI0MODE        : out std_logic;
      SPI0SSI         : in std_logic;
      SPI0SSO         : out std_logic_vector(7 downto 0);
      UART0TXD        : out std_logic;
      UART0RXD        : in std_logic;
      I2C0SDAI        : in std_logic;
      I2C0SDAO        : out std_logic;
      I2C0SCLI        : in std_logic;
      I2C0SCLO        : out std_logic;
      SPI1DO          : out std_logic;
      SPI1DOE         : out std_logic;
      SPI1DI          : in std_logic;
      SPI1CLKI        : in std_logic;
      SPI1CLKO        : out std_logic;
      SPI1MODE        : out std_logic;
      SPI1SSI         : in std_logic;
      SPI1SSO         : out std_logic_vector(7 downto 0);
      UART1TXD        : out std_logic;
      UART1RXD        : in std_logic;
      I2C1SDAI        : in std_logic;
      I2C1SDAO        : out std_logic;
      I2C1SCLI        : in std_logic;
      I2C1SCLO        : out std_logic;
      MACTXD          : out std_logic_vector(1 downto 0);
      MACRXD          : in std_logic_vector(1 downto 0);
      MACTXEN         : out std_logic;
      MACCRSDV        : in std_logic;
      MACRXER         : in std_logic;
      MACMDI          : in std_logic;
      MACMDO          : out std_logic;
      MACMDEN         : out std_logic;
      MACMDC          : out std_logic;
      EMCCLK          : out std_logic;
      EMCCLKRTN       : in std_logic;
      EMCRDB          : in std_logic_vector(15 downto 0);
      EMCAB           : out std_logic_vector(25 downto 0);
      EMCWDB          : out std_logic_vector(15 downto 0);
      EMCRWn          : out std_logic;
      EMCCS0n         : out std_logic;
      EMCCS1n         : out std_logic;
      EMCOEN0n        : out std_logic;
      EMCOEN1n        : out std_logic;
      EMCBYTEN        : out std_logic_vector(1 downto 0);
      EMCDBOE         : out std_logic;
      ADC0         : in std_logic;
      ADC1         : in std_logic;
      ADC2         : in std_logic;
      ADC3         : in std_logic;
      ADC4         : in std_logic;
      ADC5         : in std_logic;
      ADC6         : in std_logic;
      ADC7         : in std_logic;
      ADC8         : in std_logic;
      ADC9         : in std_logic;
      ADC10         : in std_logic;
      ADC11         : in std_logic;
      SDD0            : out std_logic;
      SDD1            : out std_logic;
      SDD2            : out std_logic;
      ABPS0       : in std_logic;
      ABPS1       : in std_logic;
      ABPS2       : in std_logic;
      ABPS3       : in std_logic;
      ABPS4       : in std_logic;
      ABPS5       : in std_logic;
      ABPS6       : in std_logic;
      ABPS7       : in std_logic;
      ABPS8       : in std_logic;
      ABPS9       : in std_logic;
      ABPS10       : in std_logic;
      ABPS11       : in std_logic;
      TM0          : in std_logic;
      TM1          : in std_logic;
      TM2          : in std_logic;
      TM3          : in std_logic;
      TM4          : in std_logic;
      TM5          : in std_logic;
      CM0          : in std_logic;
      CM1          : in std_logic;
      CM2          : in std_logic;
      CM3          : in std_logic;
      CM4          : in std_logic;
      CM5          : in std_logic;
      GNDTM0         : in std_logic;
      GNDTM1         : in std_logic;
      GNDTM2         : in std_logic;
      VAREF0          : in std_logic;
      VAREF1          : in std_logic;
      VAREF2          : in std_logic;
      VAREFOUT        : out std_logic;
      GNDVAREF        : in std_logic;
      PUn             : in std_logic
   );
END COMPONENT;

COMPONENT MSS_APB
  generic (
    ACT_CONFIG : integer := 0 ;
    ACT_FCLK   : integer  := 0 ;
    ACT_DIE   : string  := "" ;
    ACT_PKG   : string  := "");
   port (
      MSSPADDR        : out std_logic_vector(19 downto 0);
      MSSPWDATA       : out std_logic_vector(31 downto 0);
      MSSPWRITE       : out std_logic;
      MSSPSEL         : out std_logic;
      MSSPENABLE      : out std_logic;
      MSSPRDATA       : in std_logic_vector(31 downto 0);
      MSSPREADY       : in std_logic;
      MSSPSLVERR      : in std_logic;
      FABPADDR        : in std_logic_vector(31 downto 0);
      FABPWDATA       : in std_logic_vector(31 downto 0);
      FABPWRITE       : in std_logic;
      FABPSEL         : in std_logic;
      FABPENABLE      : in std_logic;
      FABPRDATA       : out std_logic_vector(31 downto 0);
      FABPREADY       : out std_logic;
      FABPSLVERR      : out std_logic;
      SYNCCLKFDBK     : in std_logic;
      CALIBOUT        : out std_logic;
      CALIBIN         : in std_logic;
      FABINT          : in std_logic;
      MSSINT          : out std_logic_vector(7 downto 0);
      WDINT           : out std_logic;
      F2MRESETn       : in std_logic;
      DMAREADY        : in std_logic_vector(1 downto 0);
      RXEV            : in std_logic;
      VRON            : in std_logic;
      M2FRESETn       : out std_logic;
      DEEPSLEEP       : out std_logic;
      SLEEP           : out std_logic;
      TXEV            : out std_logic;
      UART0CTSn       : in std_logic;
      UART0DSRn       : in std_logic;
      UART0RIn        : in std_logic;
      UART0DCDn       : in std_logic;
      UART0RTSn       : out std_logic;
      UART0DTRn       : out std_logic;
      UART1CTSn       : in std_logic;
      UART1DSRn       : in std_logic;
      UART1RIn        : in std_logic;
      UART1DCDn       : in std_logic;
      UART1RTSn       : out std_logic;
      UART1DTRn       : out std_logic;
      I2C0SMBUSNI     : in std_logic;
      I2C0SMBALERTNI  : in std_logic;
      I2C0BCLK        : in std_logic;
      I2C0SMBUSNO     : out std_logic;
      I2C0SMBALERTNO  : out std_logic;
      I2C1SMBUSNI     : in std_logic;
      I2C1SMBALERTNI  : in std_logic;
      I2C1BCLK        : in std_logic;
      I2C1SMBUSNO     : out std_logic;
      I2C1SMBALERTNO  : out std_logic;
      MACM2FTXD          : out std_logic_vector(1 downto 0);
      MACF2MRXD          : in std_logic_vector(1 downto 0);
      MACM2FTXEN         : out std_logic;
      MACF2MCRSDV        : in std_logic;
      MACF2MRXER         : in std_logic;
      MACF2MMDI          : in std_logic;
      MACM2FMDO          : out std_logic;
      MACM2FMDEN         : out std_logic;
      MACM2FMDC          : out std_logic;
      FABSDD0D        : in std_logic;
      FABSDD1D        : in std_logic;
      FABSDD2D        : in std_logic;
      FABSDD0CLK      : in std_logic;
      FABSDD1CLK      : in std_logic;
      FABSDD2CLK      : in std_logic;
      FABACETRIG      : in std_logic;
      ACEFLAGS  : out std_logic_vector(31 downto 0);
      CMP0            : out std_logic;
      CMP1            : out std_logic;
      CMP2            : out std_logic;
      CMP3            : out std_logic;
      CMP4            : out std_logic;
      CMP5            : out std_logic;
      CMP6            : out std_logic;
      CMP7            : out std_logic;
      CMP8            : out std_logic;
      CMP9            : out std_logic;
      CMP10           : out std_logic;
      CMP11           : out std_logic;
      LVTTL0EN      : in std_logic;
      LVTTL1EN      : in std_logic;
      LVTTL2EN      : in std_logic;
      LVTTL3EN      : in std_logic;
      LVTTL4EN      : in std_logic;
      LVTTL5EN      : in std_logic;
      LVTTL6EN      : in std_logic;
      LVTTL7EN      : in std_logic;
      LVTTL8EN      : in std_logic;
      LVTTL9EN      : in std_logic;
      LVTTL10EN     : in std_logic;
      LVTTL11EN     : in std_logic;
      LVTTL0        : out std_logic;
      LVTTL1        : out std_logic;
      LVTTL2        : out std_logic;
      LVTTL3        : out std_logic;
      LVTTL4        : out std_logic;
      LVTTL5        : out std_logic;
      LVTTL6        : out std_logic;
      LVTTL7        : out std_logic;
      LVTTL8        : out std_logic;
      LVTTL9        : out std_logic;
      LVTTL10       : out std_logic;
      LVTTL11       : out std_logic;
      PUFABn          : out std_logic;
      VCC15GOOD        : out std_logic;
      VCC33GOOD        : out std_logic;
      FCLK          : in std_logic;
      MACCLKCCC       : in std_logic;
      RCOSC           : in std_logic;
      MACCLK          : in std_logic;
      PLLLOCK         : in std_logic;
      MSSRESETn       : in std_logic;
      GPI             : in std_logic_vector(31 downto 0);
      GPO             : out std_logic_vector(31 downto 0);
      GPOE            : out std_logic_vector(31 downto 0);
      SPI0DO          : out std_logic;
      SPI0DOE         : out std_logic;
      SPI0DI          : in std_logic;
      SPI0CLKI        : in std_logic;
      SPI0CLKO        : out std_logic;
      SPI0MODE        : out std_logic;
      SPI0SSI         : in std_logic;
      SPI0SSO         : out std_logic_vector(7 downto 0);
      UART0TXD        : out std_logic;
      UART0RXD        : in std_logic;
      I2C0SDAI        : in std_logic;
      I2C0SDAO        : out std_logic;
      I2C0SCLI        : in std_logic;
      I2C0SCLO        : out std_logic;
      SPI1DO          : out std_logic;
      SPI1DOE         : out std_logic;
      SPI1DI          : in std_logic;
      SPI1CLKI        : in std_logic;
      SPI1CLKO        : out std_logic;
      SPI1MODE        : out std_logic;
      SPI1SSI         : in std_logic;
      SPI1SSO         : out std_logic_vector(7 downto 0);
      UART1TXD        : out std_logic;
      UART1RXD        : in std_logic;
      I2C1SDAI        : in std_logic;
      I2C1SDAO        : out std_logic;
      I2C1SCLI        : in std_logic;
      I2C1SCLO        : out std_logic;
      MACTXD          : out std_logic_vector(1 downto 0);
      MACRXD          : in std_logic_vector(1 downto 0);
      MACTXEN         : out std_logic;
      MACCRSDV        : in std_logic;
      MACRXER         : in std_logic;
      MACMDI          : in std_logic;
      MACMDO          : out std_logic;
      MACMDEN         : out std_logic;
      MACMDC          : out std_logic;
      EMCCLK          : out std_logic;
      EMCCLKRTN       : in std_logic;
      EMCRDB          : in std_logic_vector(15 downto 0);
      EMCAB           : out std_logic_vector(25 downto 0);
      EMCWDB          : out std_logic_vector(15 downto 0);
      EMCRWn          : out std_logic;
      EMCCS0n         : out std_logic;
      EMCCS1n         : out std_logic;
      EMCOEN0n        : out std_logic;
      EMCOEN1n        : out std_logic;
      EMCBYTEN        : out std_logic_vector(1 downto 0);
      EMCDBOE         : out std_logic;
      ADC0         : in std_logic;
      ADC1         : in std_logic;
      ADC2         : in std_logic;
      ADC3         : in std_logic;
      ADC4         : in std_logic;
      ADC5         : in std_logic;
      ADC6         : in std_logic;
      ADC7         : in std_logic;
      ADC8         : in std_logic;
      ADC9         : in std_logic;
      ADC10         : in std_logic;
      ADC11         : in std_logic;
      SDD0            : out std_logic;
      SDD1            : out std_logic;
      SDD2            : out std_logic;
      ABPS0       : in std_logic;
      ABPS1       : in std_logic;
      ABPS2       : in std_logic;
      ABPS3       : in std_logic;
      ABPS4       : in std_logic;
      ABPS5       : in std_logic;
      ABPS6       : in std_logic;
      ABPS7       : in std_logic;
      ABPS8       : in std_logic;
      ABPS9       : in std_logic;
      ABPS10       : in std_logic;
      ABPS11       : in std_logic;
      TM0          : in std_logic;
      TM1          : in std_logic;
      TM2          : in std_logic;
      TM3          : in std_logic;
      TM4          : in std_logic;
      TM5          : in std_logic;
      CM0          : in std_logic;
      CM1          : in std_logic;
      CM2          : in std_logic;
      CM3          : in std_logic;
      CM4          : in std_logic;
      CM5          : in std_logic;
      GNDTM0         : in std_logic;
      GNDTM1         : in std_logic;
      GNDTM2         : in std_logic;
      VAREF0          : in std_logic;
      VAREF1          : in std_logic;
      VAREF2          : in std_logic;
      VAREFOUT        : out std_logic;
      GNDVAREF        : in std_logic;
      PUn             : in std_logic
   );
END COMPONENT;

COMPONENT MSS_CCC
  generic (
    VCOFREQUENCY : real := 0.0 );
  port (
    CLKA         : in    std_ulogic;
    EXTFB        : in    std_ulogic;
    GLA          : out   std_ulogic;
    GLAMSS       : out   std_ulogic;
    LOCK         : out   std_ulogic;
    LOCKMSS      : out   std_ulogic;
    CLKB         : in    std_ulogic;
    GLB          : out   std_ulogic;
    YB           : out   std_ulogic;
    CLKC         : in    std_ulogic;
    GLC          : out   std_ulogic;
    YC           : out   std_ulogic;
    MACCLK       : out   std_ulogic;
    OADIV        : in    std_ulogic_vector(4 downto 0);
    OADIVHALF    : in    std_ulogic;
    OAMUX        : in    std_ulogic_vector(2 downto 0);
    BYPASSA      : in    std_ulogic;
    DLYGLA       : in    std_ulogic_vector(4 downto 0);
    DLYGLAMSS    : in    std_ulogic_vector(4 downto 0);
    DLYGLAFAB    : in    std_ulogic_vector(4 downto 0);
    OBDIV        : in    std_ulogic_vector(4 downto 0);
    OBDIVHALF    : in    std_ulogic;
    OBMUX        : in    std_ulogic_vector(2 downto 0);
    BYPASSB      : in    std_ulogic;
    DLYGLB       : in    std_ulogic_vector(4 downto 0);
    OCDIV        : in    std_ulogic_vector(4 downto 0);
    OCDIVHALF    : in    std_ulogic;
    OCMUX        : in    std_ulogic_vector(2 downto 0);
    BYPASSC      : in    std_ulogic;
    DLYGLC       : in    std_ulogic_vector(4 downto 0);
    FINDIV       : in    std_ulogic_vector(6 downto 0);
    FBDIV        : in    std_ulogic_vector(6 downto 0);
    FBDLY        : in    std_ulogic_vector(4 downto 0);
    FBSEL        : in    std_ulogic_vector(1 downto 0);
    XDLYSEL      : in    std_ulogic;
    GLMUXSEL     : in    std_ulogic_vector(1 downto 0);
    GLMUXCFG     : in    std_ulogic_vector(1 downto 0)
   );
  
END COMPONENT;

COMPONENT FAB_CCC
  generic (
    VCOFREQUENCY : real := 0.0 );

  port (
    CLKA         : in    std_ulogic;
    EXTFB        : in    std_ulogic;
    PLLEN        : in    std_ulogic;
    GLA          : out   std_ulogic;
    LOCK         : out   std_ulogic;
    CLKB         : in    std_ulogic;
    GLB          : out   std_ulogic;
    YB           : out   std_ulogic;
    CLKC         : in    std_ulogic;
    GLC          : out   std_ulogic;
    YC           : out   std_ulogic;
    OADIV        : in    std_ulogic_vector(4 downto 0);
    OADIVHALF    : in    std_ulogic;
    OADIVRST     : in    std_ulogic;
    OAMUX        : in    std_ulogic_vector(2 downto 0);
    BYPASSA      : in    std_ulogic;
    DLYGLA       : in    std_ulogic_vector(4 downto 0);
    DLYGLAFAB    : in    std_ulogic_vector(4 downto 0);
    OBDIV        : in    std_ulogic_vector(4 downto 0);
    OBDIVHALF    : in    std_ulogic;
    OBDIVRST     : in    std_ulogic;
    OBMUX        : in    std_ulogic_vector(2 downto 0);
    BYPASSB      : in    std_ulogic;
    DLYGLB       : in    std_ulogic_vector(4 downto 0);
    OCDIV        : in    std_ulogic_vector(4 downto 0);
    OCDIVHALF    : in    std_ulogic;
    OCDIVRST     : in    std_ulogic;
    OCMUX        : in    std_ulogic_vector(2 downto 0);
    BYPASSC      : in    std_ulogic;
    DLYGLC       : in    std_ulogic_vector(4 downto 0);
    FINDIV       : in    std_ulogic_vector(6 downto 0);
    FBDIV        : in    std_ulogic_vector(6 downto 0);
    FBDLY        : in    std_ulogic_vector(4 downto 0);
    FBSEL        : in    std_ulogic_vector(1 downto 0);
    XDLYSEL      : in    std_ulogic;
    VCOSEL       : in    std_ulogic_vector(2 downto 0);
    GLMUXINT     : in    std_ulogic;
    GLMUXSEL     : in    std_ulogic_vector(1 downto 0);
    GLMUXCFG     : in    std_ulogic_vector(1 downto 0)
   );
  
END COMPONENT;

COMPONENT FAB_CCC_DYN
  generic (
    VCOFREQUENCY : real := 0.0 );

  port (
    CLKA         : in    std_ulogic;
    EXTFB        : in    std_ulogic;
    PLLEN        : in    std_ulogic;
    GLA          : out   std_ulogic;
    LOCK         : out   std_ulogic;
    CLKB         : in    std_ulogic;
    GLB          : out   std_ulogic;
    YB           : out   std_ulogic;
    CLKC         : in    std_ulogic;
    GLC          : out   std_ulogic;
    YC           : out   std_ulogic;
    SDIN         : in    std_ulogic;
    SCLK         : in    std_ulogic;
    SSHIFT       : in    std_ulogic;
    SUPDATE      : in    std_ulogic;
    MODE         : in    std_ulogic;
    SDOUT        : out   std_ulogic;
    OADIV        : in    std_ulogic_vector(4 downto 0);
    OADIVHALF    : in    std_ulogic;
    OADIVRST     : in    std_ulogic;
    OAMUX        : in    std_ulogic_vector(2 downto 0);
    BYPASSA      : in    std_ulogic;
    DLYGLA       : in    std_ulogic_vector(4 downto 0);
    DLYGLAFAB    : in    std_ulogic_vector(4 downto 0);
    OBDIV        : in    std_ulogic_vector(4 downto 0);
    OBDIVHALF    : in    std_ulogic;
    OBDIVRST     : in    std_ulogic;
    OBMUX        : in    std_ulogic_vector(2 downto 0);
    BYPASSB      : in    std_ulogic;
    DLYGLB       : in    std_ulogic_vector(4 downto 0);
    OCDIV        : in    std_ulogic_vector(4 downto 0);
    OCDIVHALF    : in    std_ulogic;
    OCDIVRST     : in    std_ulogic;
    OCMUX        : in    std_ulogic_vector(2 downto 0);
    BYPASSC      : in    std_ulogic;
    DLYGLC       : in    std_ulogic_vector(4 downto 0);
    FINDIV       : in    std_ulogic_vector(6 downto 0);
    FBDIV        : in    std_ulogic_vector(6 downto 0);
    FBDLY        : in    std_ulogic_vector(4 downto 0);
    FBSEL        : in    std_ulogic_vector(1 downto 0);
    XDLYSEL      : in    std_ulogic;
    VCOSEL       : in    std_ulogic_vector(2 downto 0);
    GLMUXINT     : in    std_ulogic;
    GLMUXSEL     : in    std_ulogic_vector(1 downto 0);
    GLMUXCFG     : in    std_ulogic_vector(1 downto 0)
   );
  
END COMPONENT;


END COMPONENTS;
